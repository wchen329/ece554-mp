/* Small auto testbench for Convolution Filter
 * Conv. Filter
 */
module Convolution_Filter_tb();


	/* Execution
	 */
	initial begin
		
	end

endmodule
